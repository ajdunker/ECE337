/home/ecegrid/a/mg118/ece337/Lab2/source/adder_8bit.sv