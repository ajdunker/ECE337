// $Id: $
// File name:   flex_counter.sv
// Created:     2/4/2016
// Author:      Alexander Dunker
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Flexible and Scalable Counter with Controlled Rollover.
