// $Id: $
// File name:   rcu.sv
// Created:     2/11/2016
// Author:      Alexander Dunker
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Receiver control unit. Dictates the current mode of operation for the receiver block.
