// $Id: $
// File name:   tb_mealy.sv
// Created:     2/11/2016
// Author:      Alexander Dunker
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Test bench for Mealy Machine '1101' detector.
