// $Id: $
// File name:   flex_stp_sr.sv
// Created:     2/3/2016
// Author:      Alexander Dunker
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: N-bit Serial-to-Parallel Shift Register Design.
