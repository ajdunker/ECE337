// $Id: $
// File name:   rcv_block.sv
// Created:     2/11/2016
// Author:      Alexander Dunker
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Receiver block.

module rcv_block
  (
   input wire 	     clk;
   input wire 	     n_rst;
   input wire 	     serial_in;
   input wire 	     data_read;
   output wire [7:0] rx_data;
   output wire 	     ovverun_error;
   output wire 	     framing_error;
   );

   
   


end module
