// $Id: $
// File name:   sync_high.sv
// Created:     1/27/2016
// Author:      Alexander Dunker
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Reset to Logic High Synchronizer
