/home/ecegrid/a/mg118/ece337/Lab2/source/tb_adder_1bit.sv